.title KiCad schematic
.include "C:/AE/ZXCT1030/_models/BZX84C4V7.spice.txt"
.include "C:/AE/ZXCT1030/_models/C2012C0G2A102J060AA_p.mod"
.include "C:/AE/ZXCT1030/_models/C2012CH2A103J125AA_p.mod"
.include "C:/AE/ZXCT1030/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/ZXCT1030/_models/C3225X7S1H106M250AB_p.mod"
.include "C:/AE/ZXCT1030/_models/US1M.spice.txt"
.include "C:/AE/ZXCT1030/_models/ZXCT1030.spice.txt"
.include "C:/AE/ZXCT1030/_models/ZXMN3B14F.spice.txt"
.include "C:/AE/ZXCT1030/_models/ZXMP3A17E6.spice.txt"
R7 /VOCM /CURRENT_FEEDBACK {RLPF}
V1 /VIN 0 {VSOURCE}
XU4 /VIN /VSN C2012C0G2A102J060AA_p
XU6 VDD /VSN /VIN 0 /TRP unconnected-_U6-REF-Pad6_ /VOCM /COMP_OUT ZXCT1030
XU3 VDD 0 C2012X7R2A104K125AA_p
XU2 VDD 0 C3225X7S1H106M250AB_p
R1 /VIN /OCP {RSENSE1}
R2 /VIN /OCP {RSENSE2}
XU1 /VOUT /DRAIN /OCP ZXMP3A17E6
R3 /OCP /DRAIN {RGP}
R6 /COMP_OUT /GATE {RGN}
D1 /GATE /COMP_OUT DI_US1M
R4 /OCP /VSN {RLIM}
R5 VDD /COMP_OUT {RPU}
XU5 /DRAIN /GATE 0 ZXMN3B14F
R11 /TRP 0 {RREF}
R9 VDD /TRP {RADJ}
V2 VDD 0 {VSUPPLY}
XU7 0 /CURRENT_FEEDBACK DI_BZX84C4V7
XU8 /CURRENT_FEEDBACK 0 C2012CH2A103J125AA_p
S1 /OL /VOUT /VOL 0 SWITCH
V3 /VOL 0 PULSE(0 1 0.5m 50n 50n 1m 2m)
R12 /VOUT 0 {RLOAD}
R8 /OL 0 {ROL}
.end
