.title KiCad schematic
.include "C:/AE/ZXCT1030/_models/C2012C0G2A102J060AA_p.mod"
.include "C:/AE/ZXCT1030/_models/C2012CH2A103J125AA_p.mod"
.include "C:/AE/ZXCT1030/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/ZXCT1030/_models/C3225X7S1H106M250AB_p.mod"
.include "C:/AE/ZXCT1030/_models/ZXCT1030.spice.txt"
V1 /VIN 0 {VSOURCE}
XU2 VDD 0 C2012X7R2A104K125AA_p
R5 /CURRENT_FEEDBACK /VOCM {RLPF}
XU1 VDD 0 C3225X7S1H106M250AB_p
R1 /VIN /VOUT {RSENSE1}
R2 /VIN /VOUT {RSENSE2}
I1 /VOUT 0 {ILOAD}
R4 VDD /ALARM {RPU}
XU3 VDD /SN /VIN 0 /TRP unconnected-_U3-REF-Pad6_ /VOCM /ALARM ZXCT1030
R3 /VOUT /SN {RLIM}
XU5 /VIN /SN C2012CH2A103J125AA_p
R7 /TRP 0 {RREF}
R6 VDD /TRP {RADJ}
XU4 /CURRENT_FEEDBACK 0 C2012C0G2A102J060AA_p
V2 VDD 0 {VSUPPLY}
.end
