.title KiCad schematic
.include "models/BZX84C4V7.spice.txt"
.include "models/C2012C0G2A102J060AA_p.mod"
.include "models/C2012CH2A103J125AA_p.mod"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/C3225X7S1H106M250AB_p.mod"
.include "models/US1M.spice.txt"
.include "models/ZXCT1030.spice.txt"
.include "models/ZXMN3B14F.spice.txt"
.include "models/ZXMP3A17E6.spice.txt"
XU6 VDD /VSN /VIN 0 /TRP unconnected-_U6-Pad6_ /VOCM /COMP_OUT ZXCT1030
XU4 /VIN /VSN C2012C0G2A102J060AA_p
R4 /OCP /VSN {RLIM}
R1 /VIN /OCP {RSENSE1}
R2 /VIN /OCP {RSENSE2}
D1 /GATE /COMP_OUT DI_US1M
R3 /OCP /DRAIN {RGP}
XU1 /VOUT /DRAIN /OCP ZXMP3A17E6
R5 VDD /COMP_OUT {RPU}
R6 /COMP_OUT /GATE {RGN}
R12 /VOUT 0 {RLOAD}
XU5 /DRAIN /GATE 0 ZXMN3B14F
XU2 VDD 0 C3225X7S1H106M250AB_p
XU3 VDD 0 C2012X7R2A104K125AA_p
R7 /VOCM /CURRENT_FEEDBACK {RLPF}
V1 /VIN 0 {VSOURCE}
XU7 0 /CURRENT_FEEDBACK DI_BZX84C4V7
V2 VDD 0 {VSUPPLY}
R11 /TRP 0 {RREF}
R9 VDD /TRP {RADJ}
XU8 /CURRENT_FEEDBACK 0 C2012CH2A103J125AA_p
.end
